`ifndef DIV_BY_3_SEQ_ITEM
`define DIV_BY_3_SEQ_ITEM

class div_by_3_seq_item;

  //Input declared as random
  rand logic bit_number;
  rand logic res_n;
  
  //output signals
  logic divl;


endclass

`endif
