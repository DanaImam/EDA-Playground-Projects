`ifndef DIV_BY_3_IF
`define DIV_BY_3_IF

interface div_by_3_if (input logic clock);
  
  logic bit_number;
  logic res_n;
  logic divl;
  
endinterface

`endif
